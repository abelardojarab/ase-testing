class bogus;
endclass

